module main (nSimulacao ,cBotoes ,chaveNP, chaveTime ,clock ,buzzer ,led ,display);
	
	//Botoes de entrada
	//numeros de simulação simulação
	//somador
	//comparador de magnitude
	
	
//
	
	
	//btnsEntrada nSomar ( .A(cBotoes[0]), .B(cBotoes[1]), .C(cBotoes[2]), .N(//Colocar saida));
	//somadorSubtrator7bts somador (.A(nSimulacao), .B(//saidaBotoes), .Cin(chaveNP), .S(//saida soma), .Cout());

	
endmodule 