module decod7segs(BCD, n7Segs);
	
	input [3:0] BCD;
	output [6:0] n7Segs;
	
	//	A = 0010 + 0011 + 0101 + 0110 + 0111 + 1000 + 1001
	// B = 0001 + 0010 + 0011 + 0100 + 0111 + 1000 + 1001
	// C = 0001 + 0011 + 0100 + 0101 + 0110 + 0111 + 1000 + 1001
	// D = 0010 + 0011 + 0101 + 0110 + 1000 + 1001
	// E = 0010 + 0101 + 0110 + 1000
	// F = 0100 + 0110 + 1000 + 1001
	// G = 0010 + 0011 + 0100 + 0101 + 0110 + 1000 + 1001
	
	wire N0, N1, N2, N3;
	not (N3, BCD[3]);
	not (N2, BCD[2]);
	not (N1, BCD[1]);
	not (N0, BCD[0]);
	
	
	//	ANDS 1 A 9 EM BCD
	wire A0, A1, A2, A3, A4, A5, A6, A7, A8, A9 ;
	and ands00 (A0, N3 , N2, N1, N0);
	and ands01 (A1, N3 , N2, N1, BCD[0]);
	and ands02 (A2, N3 , N2, BCD[1], N0);
	and ands03 (A3, N3 , N2, BCD[1], BCD[0]);
	and ands04 (A4, N3 , BCD[2], N1, N0);
	and ands05 (A5, N3 , BCD[2], N1, BCD[0]);
	and ands06 (A6, N3 , BCD[2], BCD[1] ,N0);
	and ands07 (A7, N3 , BCD[2], BCD[1], BCD[0]);
	and ands08 (A8, BCD[3] , N2, N1, N0);
	and ands09 (A9, BCD[3] , N2, N1, BCD[0]);
	
	
	// A = 0010 + 0011 + 0101 + 0110 + 0111 + 1000 + 1001
	// ============================= SAIDA 0 =================================  
	wire t1;
	or ors00 (t1, A2, A3, A5, A6, A7, A8, A9);
	not not0 (n7Segs[0], t1);
	
	
	//B = 0001 + 0010 + 0011 + 0100 + 0111 + 1000 + 1001
	// ============================= SAIDA 1 =================================  
	wire t2;
	or ors01 (t2, A1, A2, A3, A4, A7, A8, A9);
	not not1 (n7Segs[1], t2);
	
	
	//C = 0001 + 0011 + 0100 + 0101 + 0110 + 0111 + 1000 + 1001
	// ============================= SAIDA 2 =================================  
	wire t3;
	or ors02 (t3, A1, A3, A4, A5, A6, A7, A8, A9);
	not not2 (n7Segs[2], t3);
	
	
	//D = 0010 + 0011 + 0101 + 0110 + 1000 + 1001
	// ============================= SAIDA 3 =================================  
	wire t4;
	or ors03 (t4, A2, A3, A5, A6, A8, A9);
	not not3 (n7Segs[3], t4);
	
	
	//E = 0010 + 0101 + 0110 + 1000
	// ============================= SAIDA 4 =================================  
	wire t5;
	or ors04 (t5, A2, A5, A6, A8);
	not not4 (n7Segs[4], t5);
	
	
	//F = 0100 + 0110 + 1000 + 1001
	// ============================= SAIDA 5 =================================  
	wire t6;
	or ors05 (t6, A4, A6, A8, A9);
	not not5 (n7Segs[5], t6);
	
	
	//G = 0010 + 0011 + 0100 + 0101 + 0110 + 1000 + 1001
	// ============================= SAIDA 6 =================================  
	wire t7;
	or ors06 (t7,A0, A2, A3, A4, A5, A6, A8, A9);
	not not6 (n7Segs[6], t7);
	
endmodule 