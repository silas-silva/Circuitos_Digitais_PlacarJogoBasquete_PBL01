module mainTeste(/*clock_in, resetNumero, chaveParar, chaveEscolherCronometro , saida, buzzer*/
	  );
	
//	input clock_in, resetNumero, chaveParar, chaveEscolherCronometro;
//	output [4:0] saida;
//	output buzzer;
	
//	cronometroRegressivoGeral(.clock_in(clock_in), .resetNumero(resetNumero), .chaveParar(chaveParar), .chaveEscolherCronometro(chaveEscolherCronometro) , .saida(saida), .buzzer(buzzer));
	
	
	
endmodule 